library verilog;
use verilog.vl_types.all;
entity lab1_vhdl2_vlg_check_tst is
    port(
        g               : in     vl_logic;
        h               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab1_vhdl2_vlg_check_tst;

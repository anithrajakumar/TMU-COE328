library verilog;
use verilog.vl_types.all;
entity lab1_vhdl2 is
    port(
        w1              : in     vl_logic;
        w2              : in     vl_logic;
        w3              : in     vl_logic;
        w4              : in     vl_logic;
        g               : out    vl_logic;
        h               : out    vl_logic
    );
end lab1_vhdl2;
